module main();
    HelloWorld helloWorld();
endmodule
