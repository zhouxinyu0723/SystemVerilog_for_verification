module helloWorld();
    initial begin
        $display("Hello World.");
        $finish;
    end
endmodule
